library verilog;
use verilog.vl_types.all;
entity sdr_test_vlg_vec_tst is
end sdr_test_vlg_vec_tst;
